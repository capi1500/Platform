ObjectNumber 1
Object{
position 0 0
}
End