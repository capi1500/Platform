Ground{
    position 110 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 210 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 170 110
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 50 150
    size 150 10
    shape box
    texture Textures/ground.png
}
Ground{
    position 200 150
    size 150 10
    shape box
    texture Textures/ground.png
}
Ground{
    position 350 150
    size 150 10
    shape box
    texture Textures/ground.png
}
Collectible{
    position 175 95
    size 10 10
    shape box
    type kinematic
    name Point
    texture Textures/yellowBox.png
}
Ground{
    position 500 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 520 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 540 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 560 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 580 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 600 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 620 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 640 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 660 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Ground{
    position 680 130
    size 20 20
    shape box
    texture Textures/redBox.png
}
Player{
    position 125 128
    size 19 19
    friction 0
    density 1
    shape circle
    name Player
    texture Textures/blueBox.png
}
Object{
    position 220 90
    size 20 20
    friction 0.3
    density 1
    shape box
    type dynamic
    texture Textures/redBox.png
}