time 0
Ground{
	type static
	shape box
	position 110 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 210 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 170 110
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 50 150
	size 150 10
	velocity 0 0
	angle 0
	texture Textures/ground.png
}
Ground{
	type static
	shape box
	position 200 150
	size 150 10
	velocity 0 0
	angle 0
	texture Textures/ground.png
}
Ground{
	type static
	shape box
	position 350 150
	size 150 10
	velocity 0 0
	angle 0
	texture Textures/ground.png
}
Collectible{
	type kinematic
	shape box
	position 175 95
	size 10 10
	velocity 0 0
	angle 0
	sound Audio/laser.ogg
	texture Textures/yellowBox.png
	collected false
}
Ground{
	type static
	shape box
	position 500 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 520 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 540 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 560 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 580 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 600 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 620 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 640 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 660 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Ground{
	type static
	shape box
	position 680 130
	size 20 20
	velocity 0 0
	angle 0
	texture Textures/redBox.png
}
Player{
	type dynamic
	density 1
	friction 0
	shape circle
	position 325.371 98.6773
	size 19 19
	velocity -100 -5.38538
	angle 0
	sound Audio/jump.ogg
	texture Textures/blueBox.png
	EQ{
		Point 0
	}
}
Object{
	type dynamic
	density 1
	friction 5
	shape box
	position 229.838 109.6
	size 20 20
	velocity 0 0
	angle 89.9996
	texture Textures/redBox.png
}
Object{
	type dynamic
	density 1
	friction 5
	shape box
	position 236.786 129.8
	size 20 20
	velocity 0 0
	angle 6.75523e-05
	texture Textures/redBox.png
}
Object{
	type dynamic
	density 1
	friction 5
	shape box
	position 313.688 129.8
	size 20 20
	velocity 0 0
	angle 89.9999
	texture Textures/redBox.png
}
Object{
	type dynamic
	density 1
	friction 5
	shape box
	position 265.364 129.8
	size 20 20
	velocity 0 0
	angle 0.00157031
	texture Textures/redBox.png
}
